library verilog;
use verilog.vl_types.all;
entity sc_computer_vlg_vec_tst is
end sc_computer_vlg_vec_tst;
